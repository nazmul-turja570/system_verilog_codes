class stimulus;

    function new();
        //$display("Inside Stimulus New function @ %0t", $time);
    endfunction

    // Stimulus Items
    rand bit value;

endclass
