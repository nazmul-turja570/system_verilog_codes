interface intf_cnt(input clock);

    // Internal wires/logics
    logic       data;
    logic       reset;
    logic [3:0] count;

endinterface
